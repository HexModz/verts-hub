getgenv().Enabled = true
getgenv().Theme = {
    ['Main-Color'] = Color3.fromRGB(17, 17, 17),
    ['Slider-Color'] = Color3.fromRGB(117, 34, 17),
    ['ZIndex'] = 2,
    ['Transparency'] = 1,
    ['webmUrl'] = 'https://cdn.discordapp.com/attachments/729443067647623219/887003883916886086/7tUwRI1Nd4txRDM.webm',
    ['Animated'] = true,
    ['Image-Size'] = UDim2.new(0, 618, 0, 291),
    ['Image-Pos'] = UDim2.new(0, 0, 0.135, 0)
}