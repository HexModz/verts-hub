{"VHID":"eat grass son","HWID":"Mum sheeesh"}
