{"VHID":"MHoGQTEkzEQHVuWm","HWID":"4f60f438e86b898f1ffba04c9ee2cec8badadb176337dbe4b12c213d82eeae3a82fa83c5c1a1ca7a72f7dd38954e849e979682ca62741696100c9bad31435742"}